(* blackbox *)
module sky130_fd_sc_hd__diode_2 (DIODE);
    input DIODE;
endmodule
