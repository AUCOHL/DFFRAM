VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM_5Kx32
  CLASS BLOCK ;
  FOREIGN RAM_5Kx32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2889.180 BY 2587.390 ;
  PIN A[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2247.380 0.000 2247.660 4.000 ;
    END
  END A[0]
  PIN A[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2596.980 0.000 2597.260 4.000 ;
    END
  END A[10]
  PIN A[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.940 0.000 2632.220 4.000 ;
    END
  END A[11]
  PIN A[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2666.900 0.000 2667.180 4.000 ;
    END
  END A[12]
  PIN A[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2282.340 0.000 2282.620 4.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2317.300 0.000 2317.580 4.000 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2352.260 0.000 2352.540 4.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2387.220 0.000 2387.500 4.000 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2422.180 0.000 2422.460 4.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2457.140 0.000 2457.420 4.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2492.100 0.000 2492.380 4.000 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2527.060 0.000 2527.340 4.000 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2562.020 0.000 2562.300 4.000 ;
    END
  END A[9]
  PIN CLK
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2701.860 0.000 2702.140 4.000 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1129.580 0.000 1129.860 4.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1478.720 0.000 1479.000 4.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1513.680 0.000 1513.960 4.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1548.640 0.000 1548.920 4.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1583.600 0.000 1583.880 4.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1618.560 0.000 1618.840 4.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1653.520 0.000 1653.800 4.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1688.480 0.000 1688.760 4.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1723.440 0.000 1723.720 4.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1758.400 0.000 1758.680 4.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1793.360 0.000 1793.640 4.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1164.540 0.000 1164.820 4.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.320 0.000 1828.600 4.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.280 0.000 1863.560 4.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1898.240 0.000 1898.520 4.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1933.200 0.000 1933.480 4.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1968.160 0.000 1968.440 4.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2003.120 0.000 2003.400 4.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2038.080 0.000 2038.360 4.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2073.040 0.000 2073.320 4.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2108.000 0.000 2108.280 4.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2142.960 0.000 2143.240 4.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1199.500 0.000 1199.780 4.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2177.920 0.000 2178.200 4.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2212.420 0.000 2212.700 4.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1234.460 0.000 1234.740 4.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.420 0.000 1269.700 4.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.380 0.000 1304.660 4.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1339.340 0.000 1339.620 4.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1374.300 0.000 1374.580 4.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1409.260 0.000 1409.540 4.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1444.220 0.000 1444.500 4.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.780 0.000 12.060 4.000 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 360.920 0.000 361.200 4.000 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.880 0.000 396.160 4.000 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.840 0.000 431.120 4.000 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 465.800 0.000 466.080 4.000 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 500.760 0.000 501.040 4.000 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 535.720 0.000 536.000 4.000 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 570.680 0.000 570.960 4.000 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 605.640 0.000 605.920 4.000 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 640.600 0.000 640.880 4.000 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 675.560 0.000 675.840 4.000 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.280 0.000 46.560 4.000 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.520 0.000 710.800 4.000 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 745.020 0.000 745.300 4.000 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 779.980 0.000 780.260 4.000 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 814.940 0.000 815.220 4.000 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 849.900 0.000 850.180 4.000 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 884.860 0.000 885.140 4.000 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 919.820 0.000 920.100 4.000 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 954.780 0.000 955.060 4.000 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 989.740 0.000 990.020 4.000 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1024.700 0.000 1024.980 4.000 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.240 0.000 81.520 4.000 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1059.660 0.000 1059.940 4.000 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.620 0.000 1094.900 4.000 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.200 0.000 116.480 4.000 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 151.160 0.000 151.440 4.000 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 186.120 0.000 186.400 4.000 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 221.080 0.000 221.360 4.000 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 256.040 0.000 256.320 4.000 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 291.000 0.000 291.280 4.000 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 325.960 0.000 326.240 4.000 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2876.660 0.000 2876.940 4.000 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2736.820 0.000 2737.100 4.000 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2771.780 0.000 2772.060 4.000 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2806.740 0.000 2807.020 4.000 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2841.700 0.000 2841.980 4.000 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.710 10.640 17.310 2586.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 92.510 10.640 94.110 2586.960 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.190 7.225 2888.990 2586.805 ;
      LAYER met1 ;
        RECT 0.190 4.460 2888.990 2587.360 ;
      LAYER met2 ;
        RECT 1.670 4.280 2887.510 2587.390 ;
        RECT 1.670 4.000 11.500 4.280 ;
        RECT 12.340 4.000 46.000 4.280 ;
        RECT 46.840 4.000 80.960 4.280 ;
        RECT 81.800 4.000 115.920 4.280 ;
        RECT 116.760 4.000 150.880 4.280 ;
        RECT 151.720 4.000 185.840 4.280 ;
        RECT 186.680 4.000 220.800 4.280 ;
        RECT 221.640 4.000 255.760 4.280 ;
        RECT 256.600 4.000 290.720 4.280 ;
        RECT 291.560 4.000 325.680 4.280 ;
        RECT 326.520 4.000 360.640 4.280 ;
        RECT 361.480 4.000 395.600 4.280 ;
        RECT 396.440 4.000 430.560 4.280 ;
        RECT 431.400 4.000 465.520 4.280 ;
        RECT 466.360 4.000 500.480 4.280 ;
        RECT 501.320 4.000 535.440 4.280 ;
        RECT 536.280 4.000 570.400 4.280 ;
        RECT 571.240 4.000 605.360 4.280 ;
        RECT 606.200 4.000 640.320 4.280 ;
        RECT 641.160 4.000 675.280 4.280 ;
        RECT 676.120 4.000 710.240 4.280 ;
        RECT 711.080 4.000 744.740 4.280 ;
        RECT 745.580 4.000 779.700 4.280 ;
        RECT 780.540 4.000 814.660 4.280 ;
        RECT 815.500 4.000 849.620 4.280 ;
        RECT 850.460 4.000 884.580 4.280 ;
        RECT 885.420 4.000 919.540 4.280 ;
        RECT 920.380 4.000 954.500 4.280 ;
        RECT 955.340 4.000 989.460 4.280 ;
        RECT 990.300 4.000 1024.420 4.280 ;
        RECT 1025.260 4.000 1059.380 4.280 ;
        RECT 1060.220 4.000 1094.340 4.280 ;
        RECT 1095.180 4.000 1129.300 4.280 ;
        RECT 1130.140 4.000 1164.260 4.280 ;
        RECT 1165.100 4.000 1199.220 4.280 ;
        RECT 1200.060 4.000 1234.180 4.280 ;
        RECT 1235.020 4.000 1269.140 4.280 ;
        RECT 1269.980 4.000 1304.100 4.280 ;
        RECT 1304.940 4.000 1339.060 4.280 ;
        RECT 1339.900 4.000 1374.020 4.280 ;
        RECT 1374.860 4.000 1408.980 4.280 ;
        RECT 1409.820 4.000 1443.940 4.280 ;
        RECT 1444.780 4.000 1478.440 4.280 ;
        RECT 1479.280 4.000 1513.400 4.280 ;
        RECT 1514.240 4.000 1548.360 4.280 ;
        RECT 1549.200 4.000 1583.320 4.280 ;
        RECT 1584.160 4.000 1618.280 4.280 ;
        RECT 1619.120 4.000 1653.240 4.280 ;
        RECT 1654.080 4.000 1688.200 4.280 ;
        RECT 1689.040 4.000 1723.160 4.280 ;
        RECT 1724.000 4.000 1758.120 4.280 ;
        RECT 1758.960 4.000 1793.080 4.280 ;
        RECT 1793.920 4.000 1828.040 4.280 ;
        RECT 1828.880 4.000 1863.000 4.280 ;
        RECT 1863.840 4.000 1897.960 4.280 ;
        RECT 1898.800 4.000 1932.920 4.280 ;
        RECT 1933.760 4.000 1967.880 4.280 ;
        RECT 1968.720 4.000 2002.840 4.280 ;
        RECT 2003.680 4.000 2037.800 4.280 ;
        RECT 2038.640 4.000 2072.760 4.280 ;
        RECT 2073.600 4.000 2107.720 4.280 ;
        RECT 2108.560 4.000 2142.680 4.280 ;
        RECT 2143.520 4.000 2177.640 4.280 ;
        RECT 2178.480 4.000 2212.140 4.280 ;
        RECT 2212.980 4.000 2247.100 4.280 ;
        RECT 2247.940 4.000 2282.060 4.280 ;
        RECT 2282.900 4.000 2317.020 4.280 ;
        RECT 2317.860 4.000 2351.980 4.280 ;
        RECT 2352.820 4.000 2386.940 4.280 ;
        RECT 2387.780 4.000 2421.900 4.280 ;
        RECT 2422.740 4.000 2456.860 4.280 ;
        RECT 2457.700 4.000 2491.820 4.280 ;
        RECT 2492.660 4.000 2526.780 4.280 ;
        RECT 2527.620 4.000 2561.740 4.280 ;
        RECT 2562.580 4.000 2596.700 4.280 ;
        RECT 2597.540 4.000 2631.660 4.280 ;
        RECT 2632.500 4.000 2666.620 4.280 ;
        RECT 2667.460 4.000 2701.580 4.280 ;
        RECT 2702.420 4.000 2736.540 4.280 ;
        RECT 2737.380 4.000 2771.500 4.280 ;
        RECT 2772.340 4.000 2806.460 4.280 ;
        RECT 2807.300 4.000 2841.420 4.280 ;
        RECT 2842.260 4.000 2876.380 4.280 ;
        RECT 2877.220 4.000 2887.510 4.280 ;
      LAYER met3 ;
        RECT 3.015 4.255 2887.085 2586.885 ;
      LAYER met4 ;
        RECT 17.965 10.240 92.110 2586.960 ;
        RECT 94.510 10.240 2860.175 2586.960 ;
        RECT 17.965 8.335 2860.175 10.240 ;
      LAYER met5 ;
        RECT 1187.570 317.100 1813.850 2168.300 ;
  END
END RAM_5Kx32
END LIBRARY

