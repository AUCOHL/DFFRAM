VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM_4Kx32
  CLASS BLOCK ;
  FOREIGN RAM_4Kx32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2489.625 BY 2586.960 ;
  PIN A[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1960.800 0.000 1961.080 4.000 ;
    END
  END A[0]
  PIN A[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2265.780 0.000 2266.060 4.000 ;
    END
  END A[10]
  PIN A[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2296.600 0.000 2296.880 4.000 ;
    END
  END A[11]
  PIN A[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1991.620 0.000 1991.900 4.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2021.980 0.000 2022.260 4.000 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2052.340 0.000 2052.620 4.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2083.160 0.000 2083.440 4.000 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.520 0.000 2113.800 4.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.880 0.000 2144.160 4.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2174.240 0.000 2174.520 4.000 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2205.060 0.000 2205.340 4.000 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2235.420 0.000 2235.700 4.000 ;
    END
  END A[9]
  PIN CLK
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2326.960 0.000 2327.240 4.000 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 985.140 0.000 985.420 4.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1290.120 0.000 1290.400 4.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1320.940 0.000 1321.220 4.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1351.300 0.000 1351.580 4.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1381.660 0.000 1381.940 4.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.020 0.000 1412.300 4.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1442.840 0.000 1443.120 4.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1473.200 0.000 1473.480 4.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1503.560 0.000 1503.840 4.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1534.380 0.000 1534.660 4.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1564.740 0.000 1565.020 4.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1015.960 0.000 1016.240 4.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1595.100 0.000 1595.380 4.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1625.460 0.000 1625.740 4.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1656.280 0.000 1656.560 4.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1686.640 0.000 1686.920 4.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1717.000 0.000 1717.280 4.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1747.360 0.000 1747.640 4.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1778.180 0.000 1778.460 4.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1808.540 0.000 1808.820 4.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1838.900 0.000 1839.180 4.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1869.720 0.000 1870.000 4.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1046.320 0.000 1046.600 4.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1900.080 0.000 1900.360 4.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1930.440 0.000 1930.720 4.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1076.680 0.000 1076.960 4.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1107.500 0.000 1107.780 4.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1137.860 0.000 1138.140 4.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.220 0.000 1168.500 4.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1198.580 0.000 1198.860 4.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1229.400 0.000 1229.680 4.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1259.760 0.000 1260.040 4.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 9.940 0.000 10.220 4.000 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 314.460 0.000 314.740 4.000 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 345.280 0.000 345.560 4.000 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 375.640 0.000 375.920 4.000 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 406.000 0.000 406.280 4.000 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 436.360 0.000 436.640 4.000 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 467.180 0.000 467.460 4.000 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 497.540 0.000 497.820 4.000 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 527.900 0.000 528.180 4.000 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 558.720 0.000 559.000 4.000 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 589.080 0.000 589.360 4.000 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.300 0.000 40.580 4.000 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 619.440 0.000 619.720 4.000 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 649.800 0.000 650.080 4.000 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 680.620 0.000 680.900 4.000 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.980 0.000 711.260 4.000 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 741.340 0.000 741.620 4.000 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 772.160 0.000 772.440 4.000 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 802.520 0.000 802.800 4.000 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 832.880 0.000 833.160 4.000 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 863.240 0.000 863.520 4.000 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 894.060 0.000 894.340 4.000 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.660 0.000 70.940 4.000 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.420 0.000 924.700 4.000 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 954.780 0.000 955.060 4.000 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.020 0.000 101.300 4.000 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.840 0.000 132.120 4.000 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.200 0.000 162.480 4.000 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 192.560 0.000 192.840 4.000 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.920 0.000 223.200 4.000 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 253.740 0.000 254.020 4.000 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 284.100 0.000 284.380 4.000 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2479.220 0.000 2479.500 4.000 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.320 0.000 2357.600 4.000 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2387.680 0.000 2387.960 4.000 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2418.500 0.000 2418.780 4.000 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2448.860 0.000 2449.140 4.000 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.710 10.640 17.310 2586.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 92.510 10.640 94.110 2586.960 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.190 10.795 2489.565 2586.805 ;
      LAYER met1 ;
        RECT 0.190 4.800 2489.625 2586.960 ;
      LAYER met2 ;
        RECT 1.210 4.280 2487.320 2586.960 ;
        RECT 1.210 4.000 9.660 4.280 ;
        RECT 10.500 4.000 40.020 4.280 ;
        RECT 40.860 4.000 70.380 4.280 ;
        RECT 71.220 4.000 100.740 4.280 ;
        RECT 101.580 4.000 131.560 4.280 ;
        RECT 132.400 4.000 161.920 4.280 ;
        RECT 162.760 4.000 192.280 4.280 ;
        RECT 193.120 4.000 222.640 4.280 ;
        RECT 223.480 4.000 253.460 4.280 ;
        RECT 254.300 4.000 283.820 4.280 ;
        RECT 284.660 4.000 314.180 4.280 ;
        RECT 315.020 4.000 345.000 4.280 ;
        RECT 345.840 4.000 375.360 4.280 ;
        RECT 376.200 4.000 405.720 4.280 ;
        RECT 406.560 4.000 436.080 4.280 ;
        RECT 436.920 4.000 466.900 4.280 ;
        RECT 467.740 4.000 497.260 4.280 ;
        RECT 498.100 4.000 527.620 4.280 ;
        RECT 528.460 4.000 558.440 4.280 ;
        RECT 559.280 4.000 588.800 4.280 ;
        RECT 589.640 4.000 619.160 4.280 ;
        RECT 620.000 4.000 649.520 4.280 ;
        RECT 650.360 4.000 680.340 4.280 ;
        RECT 681.180 4.000 710.700 4.280 ;
        RECT 711.540 4.000 741.060 4.280 ;
        RECT 741.900 4.000 771.880 4.280 ;
        RECT 772.720 4.000 802.240 4.280 ;
        RECT 803.080 4.000 832.600 4.280 ;
        RECT 833.440 4.000 862.960 4.280 ;
        RECT 863.800 4.000 893.780 4.280 ;
        RECT 894.620 4.000 924.140 4.280 ;
        RECT 924.980 4.000 954.500 4.280 ;
        RECT 955.340 4.000 984.860 4.280 ;
        RECT 985.700 4.000 1015.680 4.280 ;
        RECT 1016.520 4.000 1046.040 4.280 ;
        RECT 1046.880 4.000 1076.400 4.280 ;
        RECT 1077.240 4.000 1107.220 4.280 ;
        RECT 1108.060 4.000 1137.580 4.280 ;
        RECT 1138.420 4.000 1167.940 4.280 ;
        RECT 1168.780 4.000 1198.300 4.280 ;
        RECT 1199.140 4.000 1229.120 4.280 ;
        RECT 1229.960 4.000 1259.480 4.280 ;
        RECT 1260.320 4.000 1289.840 4.280 ;
        RECT 1290.680 4.000 1320.660 4.280 ;
        RECT 1321.500 4.000 1351.020 4.280 ;
        RECT 1351.860 4.000 1381.380 4.280 ;
        RECT 1382.220 4.000 1411.740 4.280 ;
        RECT 1412.580 4.000 1442.560 4.280 ;
        RECT 1443.400 4.000 1472.920 4.280 ;
        RECT 1473.760 4.000 1503.280 4.280 ;
        RECT 1504.120 4.000 1534.100 4.280 ;
        RECT 1534.940 4.000 1564.460 4.280 ;
        RECT 1565.300 4.000 1594.820 4.280 ;
        RECT 1595.660 4.000 1625.180 4.280 ;
        RECT 1626.020 4.000 1656.000 4.280 ;
        RECT 1656.840 4.000 1686.360 4.280 ;
        RECT 1687.200 4.000 1716.720 4.280 ;
        RECT 1717.560 4.000 1747.080 4.280 ;
        RECT 1747.920 4.000 1777.900 4.280 ;
        RECT 1778.740 4.000 1808.260 4.280 ;
        RECT 1809.100 4.000 1838.620 4.280 ;
        RECT 1839.460 4.000 1869.440 4.280 ;
        RECT 1870.280 4.000 1899.800 4.280 ;
        RECT 1900.640 4.000 1930.160 4.280 ;
        RECT 1931.000 4.000 1960.520 4.280 ;
        RECT 1961.360 4.000 1991.340 4.280 ;
        RECT 1992.180 4.000 2021.700 4.280 ;
        RECT 2022.540 4.000 2052.060 4.280 ;
        RECT 2052.900 4.000 2082.880 4.280 ;
        RECT 2083.720 4.000 2113.240 4.280 ;
        RECT 2114.080 4.000 2143.600 4.280 ;
        RECT 2144.440 4.000 2173.960 4.280 ;
        RECT 2174.800 4.000 2204.780 4.280 ;
        RECT 2205.620 4.000 2235.140 4.280 ;
        RECT 2235.980 4.000 2265.500 4.280 ;
        RECT 2266.340 4.000 2296.320 4.280 ;
        RECT 2297.160 4.000 2326.680 4.280 ;
        RECT 2327.520 4.000 2357.040 4.280 ;
        RECT 2357.880 4.000 2387.400 4.280 ;
        RECT 2388.240 4.000 2418.220 4.280 ;
        RECT 2419.060 4.000 2448.580 4.280 ;
        RECT 2449.420 4.000 2478.940 4.280 ;
        RECT 2479.780 4.000 2487.320 4.280 ;
      LAYER met3 ;
        RECT 2.555 4.255 2487.345 2586.885 ;
      LAYER met4 ;
        RECT 9.685 10.640 15.310 2586.960 ;
        RECT 17.710 10.640 92.110 2586.960 ;
        RECT 94.510 10.640 2474.910 2586.960 ;
  END
END RAM_4Kx32
END LIBRARY

